{
  "name": "node-tachyon",
  "version": "2.1.4",
  "lockfileVersion": 1,
  "requires": true,
  "dependencies": {
    "animated-gif-detector": {
      "version": "1.2.0",
      "resolved": "https://registry.npmjs.org/animated-gif-detector/-/animated-gif-detector-1.2.0.tgz",
      "integrity": "sha1-yy+ZEcqAJPKzTGk7f9ZFQu5BYYk=",
      "requires": {
        "inherits": "2.0.3"
      }
    },
    "aws-sdk": {
      "version": "2.269.1",
      "resolved": "https://registry.npmjs.org/aws-sdk/-/aws-sdk-2.269.1.tgz",
      "integrity": "sha512-oIKzffzGR8fA9uT181wyahXQK5yBqF+qzql+0XoFePcFo7l8m8L9MAq5J9QSFXRNFM8cThjnSQpFoesVNzh7Pg==",
      "dev": true,
      "requires": {
        "buffer": "4.9.1",
        "events": "1.1.1",
        "ieee754": "1.1.8",
        "jmespath": "0.15.0",
        "querystring": "0.2.0",
        "sax": "1.2.1",
        "url": "0.10.3",
        "uuid": "3.1.0",
        "xml2js": "0.4.17"
      }
    },
    "balanced-match": {
      "version": "1.0.0",
      "resolved": "https://registry.npmjs.org/balanced-match/-/balanced-match-1.0.0.tgz",
      "integrity": "sha1-ibTRmasr7kneFk6gK4nORi1xt2c="
    },
    "base64-js": {
      "version": "1.3.0",
      "resolved": "https://registry.npmjs.org/base64-js/-/base64-js-1.3.0.tgz",
      "integrity": "sha512-ccav/yGvoa80BQDljCxsmmQ3Xvx60/UpBIij5QN21W3wBi/hhIC9OoO+KLpu9IJTS9j4DRVJ3aDDF9cMSoa2lw==",
      "dev": true
    },
    "block-stream": {
      "version": "0.0.9",
      "resolved": "https://registry.npmjs.org/block-stream/-/block-stream-0.0.9.tgz",
      "integrity": "sha1-E+v+d4oDIFz+A3UUgeu0szAMEmo=",
      "requires": {
        "inherits": "2.0.3"
      }
    },
    "brace-expansion": {
      "version": "1.1.11",
      "resolved": "https://registry.npmjs.org/brace-expansion/-/brace-expansion-1.1.11.tgz",
      "integrity": "sha512-iCuPHDFgrHX7H2vEI/5xpz07zSHB00TpugqhmYtVmMO6518mCuRMoOYFldEBl0g187ufozdaHgWKcYFb61qGiA==",
      "requires": {
        "balanced-match": "1.0.0",
        "concat-map": "0.0.1"
      }
    },
    "buffer": {
      "version": "4.9.1",
      "resolved": "https://registry.npmjs.org/buffer/-/buffer-4.9.1.tgz",
      "integrity": "sha1-bRu2AbB6TvztlwlBMgkwJ8lbwpg=",
      "dev": true,
      "requires": {
        "base64-js": "1.3.0",
        "ieee754": "1.1.8",
        "isarray": "1.0.0"
      }
    },
    "capture-stack-trace": {
      "version": "1.0.0",
      "resolved": "https://registry.npmjs.org/capture-stack-trace/-/capture-stack-trace-1.0.0.tgz",
      "integrity": "sha1-Sm+gc5nCa7pH8LJJa00PtAjFVQ0="
    },
    "caw": {
      "version": "2.0.1",
      "resolved": "https://registry.npmjs.org/caw/-/caw-2.0.1.tgz",
      "integrity": "sha512-Cg8/ZSBEa8ZVY9HspcGUYaK63d/bN7rqS3CYCzEGUxuYv6UlmcjzDUz2fCFFHyTvUW5Pk0I+3hkA3iXlIj6guA==",
      "requires": {
        "get-proxy": "2.1.0",
        "isurl": "1.0.0",
        "tunnel-agent": "0.6.0",
        "url-to-options": "1.0.1"
      }
    },
    "cli-table": {
      "version": "0.3.1",
      "resolved": "https://registry.npmjs.org/cli-table/-/cli-table-0.3.1.tgz",
      "integrity": "sha1-9TsFJmqLGguTSz0IIebi3FkUriM=",
      "dev": true,
      "requires": {
        "colors": "1.0.3"
      }
    },
    "color": {
      "version": "1.0.3",
      "resolved": "https://registry.npmjs.org/color/-/color-1.0.3.tgz",
      "integrity": "sha1-5I6DLYXxTvaU+0aIEcLVz+cptV0=",
      "requires": {
        "color-convert": "1.9.2",
        "color-string": "1.5.2"
      }
    },
    "color-convert": {
      "version": "1.9.2",
      "resolved": "https://registry.npmjs.org/color-convert/-/color-convert-1.9.2.tgz",
      "integrity": "sha512-3NUJZdhMhcdPn8vJ9v2UQJoH0qqoGUkYTgFEPZaPjEtwmmKUfNV46zZmgB2M5M4DCEQHMaCfWHCxiBflLm04Tg==",
      "requires": {
        "color-name": "1.1.1"
      }
    },
    "color-name": {
      "version": "1.1.1",
      "resolved": "https://registry.npmjs.org/color-name/-/color-name-1.1.1.tgz",
      "integrity": "sha1-SxQVMEz1ACjqgWQ2Q72C6gWANok="
    },
    "color-string": {
      "version": "1.5.2",
      "resolved": "https://registry.npmjs.org/color-string/-/color-string-1.5.2.tgz",
      "integrity": "sha1-JuRYFLw8mny9Z1FkikFDRRSnc6k=",
      "requires": {
        "color-name": "1.1.1",
        "simple-swizzle": "0.2.2"
      }
    },
    "colors": {
      "version": "1.0.3",
      "resolved": "https://registry.npmjs.org/colors/-/colors-1.0.3.tgz",
      "integrity": "sha1-BDP0TYCWgP3rYO0mDxsMJi6CpAs=",
      "dev": true
    },
    "concat-map": {
      "version": "0.0.1",
      "resolved": "https://registry.npmjs.org/concat-map/-/concat-map-0.0.1.tgz",
      "integrity": "sha1-2Klr13/Wjfd5OnMDajug1UBdR3s="
    },
    "config-chain": {
      "version": "1.1.11",
      "resolved": "https://registry.npmjs.org/config-chain/-/config-chain-1.1.11.tgz",
      "integrity": "sha1-q6CXR9++TD5w52am5BWG4YWfxvI=",
      "requires": {
        "ini": "1.3.5",
        "proto-list": "1.2.4"
      }
    },
    "create-error-class": {
      "version": "3.0.2",
      "resolved": "https://registry.npmjs.org/create-error-class/-/create-error-class-3.0.2.tgz",
      "integrity": "sha1-Br56vvlHo/FKMP1hBnHUAbyot7Y=",
      "requires": {
        "capture-stack-trace": "1.0.0"
      }
    },
    "duplexer3": {
      "version": "0.1.4",
      "resolved": "https://registry.npmjs.org/duplexer3/-/duplexer3-0.1.4.tgz",
      "integrity": "sha1-7gHdHKwO08vH/b6jfcCo8c4ALOI="
    },
    "events": {
      "version": "1.1.1",
      "resolved": "https://registry.npmjs.org/events/-/events-1.1.1.tgz",
      "integrity": "sha1-nr23Y1rQmccNzEwqH1AEKI6L2SQ=",
      "dev": true
    },
    "filesize": {
      "version": "3.6.1",
      "resolved": "https://registry.npmjs.org/filesize/-/filesize-3.6.1.tgz",
      "integrity": "sha512-7KjR1vv6qnicaPMi1iiTcI85CyYwRO/PSFCu6SvqL8jN2Wjt/NIYQTFtFs7fSDCYOstUkEWIQGFUg5YZQfjlcg==",
      "dev": true
    },
    "fs.realpath": {
      "version": "1.0.0",
      "resolved": "https://registry.npmjs.org/fs.realpath/-/fs.realpath-1.0.0.tgz",
      "integrity": "sha1-FQStJSMVjKpA20onh8sBQRmU6k8="
    },
    "fstream": {
      "version": "1.0.11",
      "resolved": "https://registry.npmjs.org/fstream/-/fstream-1.0.11.tgz",
      "integrity": "sha1-XB+x8RdHcRTwYyoOtLcbPLD9MXE=",
      "requires": {
        "graceful-fs": "4.1.11",
        "inherits": "2.0.3",
        "mkdirp": "0.5.1",
        "rimraf": "2.6.2"
      }
    },
    "get-proxy": {
      "version": "2.1.0",
      "resolved": "https://registry.npmjs.org/get-proxy/-/get-proxy-2.1.0.tgz",
      "integrity": "sha512-zmZIaQTWnNQb4R4fJUEp/FC51eZsc6EkErspy3xtIYStaq8EB/hDIWipxsal+E8rz0qD7f2sL/NA9Xee4RInJw==",
      "requires": {
        "npm-conf": "1.1.3"
      }
    },
    "get-stream": {
      "version": "3.0.0",
      "resolved": "https://registry.npmjs.org/get-stream/-/get-stream-3.0.0.tgz",
      "integrity": "sha1-jpQ9E1jcN1VQVOy+LtsFqhdO3hQ="
    },
    "glob": {
      "version": "7.1.2",
      "resolved": "https://registry.npmjs.org/glob/-/glob-7.1.2.tgz",
      "integrity": "sha512-MJTUg1kjuLeQCJ+ccE4Vpa6kKVXkPYJ2mOCQyUuKLcLQsdrMCpBPUi8qVE6+YuaJkozeA9NusTAw3hLr8Xe5EQ==",
      "requires": {
        "fs.realpath": "1.0.0",
        "inflight": "1.0.6",
        "inherits": "2.0.3",
        "minimatch": "3.0.4",
        "once": "1.4.0",
        "path-is-absolute": "1.0.1"
      }
    },
    "got": {
      "version": "6.7.1",
      "resolved": "https://registry.npmjs.org/got/-/got-6.7.1.tgz",
      "integrity": "sha1-JAzQV4WpoY5WHcG0S0HHY+8ejbA=",
      "requires": {
        "create-error-class": "3.0.2",
        "duplexer3": "0.1.4",
        "get-stream": "3.0.0",
        "is-redirect": "1.0.0",
        "is-retry-allowed": "1.1.0",
        "is-stream": "1.1.0",
        "lowercase-keys": "1.0.1",
        "safe-buffer": "5.1.2",
        "timed-out": "4.0.1",
        "unzip-response": "2.0.1",
        "url-parse-lax": "1.0.0"
      }
    },
    "graceful-fs": {
      "version": "4.1.11",
      "resolved": "https://registry.npmjs.org/graceful-fs/-/graceful-fs-4.1.11.tgz",
      "integrity": "sha1-Dovf5NHduIVNZOBOp8AOKgJuVlg="
    },
    "has-symbol-support-x": {
      "version": "1.4.2",
      "resolved": "https://registry.npmjs.org/has-symbol-support-x/-/has-symbol-support-x-1.4.2.tgz",
      "integrity": "sha512-3ToOva++HaW+eCpgqZrCfN51IPB+7bJNVT6CUATzueB5Heb8o6Nam0V3HG5dlDvZU1Gn5QLcbahiKw/XVk5JJw=="
    },
    "has-to-string-tag-x": {
      "version": "1.4.1",
      "resolved": "https://registry.npmjs.org/has-to-string-tag-x/-/has-to-string-tag-x-1.4.1.tgz",
      "integrity": "sha512-vdbKfmw+3LoOYVr+mtxHaX5a96+0f3DljYd8JOqvOLsf5mw2Otda2qCDT9qRqLAhrjyQ0h7ual5nOiASpsGNFw==",
      "requires": {
        "has-symbol-support-x": "1.4.2"
      }
    },
    "ieee754": {
      "version": "1.1.8",
      "resolved": "https://registry.npmjs.org/ieee754/-/ieee754-1.1.8.tgz",
      "integrity": "sha1-vjPUCsEO8ZJnAfbwii2G+/0a0+Q=",
      "dev": true
    },
    "inflight": {
      "version": "1.0.6",
      "resolved": "https://registry.npmjs.org/inflight/-/inflight-1.0.6.tgz",
      "integrity": "sha1-Sb1jMdfQLQwJvJEKEHW6gWW1bfk=",
      "requires": {
        "once": "1.4.0",
        "wrappy": "1.0.2"
      }
    },
    "inherits": {
      "version": "2.0.3",
      "resolved": "https://registry.npmjs.org/inherits/-/inherits-2.0.3.tgz",
      "integrity": "sha1-Yzwsg+PaQqUC9SRmAiSA9CCCYd4="
    },
    "ini": {
      "version": "1.3.5",
      "resolved": "https://registry.npmjs.org/ini/-/ini-1.3.5.tgz",
      "integrity": "sha512-RZY5huIKCMRWDUqZlEi72f/lmXKMvuszcMBduliQ3nnWbx9X/ZBQO7DijMEYS9EhHBb2qacRUMtC7svLwe0lcw=="
    },
    "is-arrayish": {
      "version": "0.3.2",
      "resolved": "https://registry.npmjs.org/is-arrayish/-/is-arrayish-0.3.2.tgz",
      "integrity": "sha512-eVRqCvVlZbuw3GrM63ovNSNAeA1K16kaR/LRY/92w0zxQ5/1YzwblUX652i4Xs9RwAGjW9d9y6X88t8OaAJfWQ=="
    },
    "is-object": {
      "version": "1.0.1",
      "resolved": "https://registry.npmjs.org/is-object/-/is-object-1.0.1.tgz",
      "integrity": "sha1-iVJojF7C/9awPsyF52ngKQMINHA="
    },
    "is-redirect": {
      "version": "1.0.0",
      "resolved": "https://registry.npmjs.org/is-redirect/-/is-redirect-1.0.0.tgz",
      "integrity": "sha1-HQPd7VO9jbDzDCbk+V02/HyH3CQ="
    },
    "is-retry-allowed": {
      "version": "1.1.0",
      "resolved": "https://registry.npmjs.org/is-retry-allowed/-/is-retry-allowed-1.1.0.tgz",
      "integrity": "sha1-EaBgVotnM5REAz0BJaYaINVk+zQ="
    },
    "is-stream": {
      "version": "1.1.0",
      "resolved": "https://registry.npmjs.org/is-stream/-/is-stream-1.1.0.tgz",
      "integrity": "sha1-EtSj3U5o4Lec6428hBc66A2RykQ="
    },
    "isarray": {
      "version": "1.0.0",
      "resolved": "https://registry.npmjs.org/isarray/-/isarray-1.0.0.tgz",
      "integrity": "sha1-u5NdSFgsuhaMBoNJV6VKPgcSTxE=",
      "dev": true
    },
    "isurl": {
      "version": "1.0.0",
      "resolved": "https://registry.npmjs.org/isurl/-/isurl-1.0.0.tgz",
      "integrity": "sha512-1P/yWsxPlDtn7QeRD+ULKQPaIaN6yF368GZ2vDfv0AL0NwpStafjWCDDdn0k8wgFMWpVAqG7oJhxHnlud42i9w==",
      "requires": {
        "has-to-string-tag-x": "1.4.1",
        "is-object": "1.0.1"
      }
    },
    "jmespath": {
      "version": "0.15.0",
      "resolved": "https://registry.npmjs.org/jmespath/-/jmespath-0.15.0.tgz",
      "integrity": "sha1-o/Iiqarp+Wb10nx5ZRDigJF2Qhc=",
      "dev": true
    },
    "lodash": {
      "version": "4.17.10",
      "resolved": "https://registry.npmjs.org/lodash/-/lodash-4.17.10.tgz",
      "integrity": "sha512-UejweD1pDoXu+AD825lWwp4ZGtSwgnpZxb3JDViD7StjQz+Nb/6l093lx4OQ0foGWNRoc19mWy7BzL+UAK2iVg==",
      "dev": true
    },
    "lowercase-keys": {
      "version": "1.0.1",
      "resolved": "https://registry.npmjs.org/lowercase-keys/-/lowercase-keys-1.0.1.tgz",
      "integrity": "sha512-G2Lj61tXDnVFFOi8VZds+SoQjtQC3dgokKdDG2mTm1tx4m50NUHBOZSBwQQHyy0V12A0JTG4icfZQH+xPyh8VA=="
    },
    "minimatch": {
      "version": "3.0.4",
      "resolved": "https://registry.npmjs.org/minimatch/-/minimatch-3.0.4.tgz",
      "integrity": "sha512-yJHVQEhyqPLUTgt9B83PXu6W3rx4MvvHvSUvToogpwoGDOUQ+yDrR0HRot+yOCdCO7u4hX3pWft6kWBBcqh0UA==",
      "requires": {
        "brace-expansion": "1.1.11"
      }
    },
    "minimist": {
      "version": "0.0.8",
      "resolved": "https://registry.npmjs.org/minimist/-/minimist-0.0.8.tgz",
      "integrity": "sha1-hX/Kv8M5fSYluCKCYuhqp6ARsF0="
    },
    "mkdirp": {
      "version": "0.5.1",
      "resolved": "https://registry.npmjs.org/mkdirp/-/mkdirp-0.5.1.tgz",
      "integrity": "sha1-MAV0OOrGz3+MR2fzhkjWaX11yQM=",
      "requires": {
        "minimist": "0.0.8"
      }
    },
    "nan": {
      "version": "2.10.0",
      "resolved": "https://registry.npmjs.org/nan/-/nan-2.10.0.tgz",
      "integrity": "sha512-bAdJv7fBLhWC+/Bls0Oza+mvTaNQtP+1RyhhhvD95pgUJz6XM5IzgmxOkItJ9tkoCiplvAnXI1tNmmUD/eScyA=="
    },
    "npm-conf": {
      "version": "1.1.3",
      "resolved": "https://registry.npmjs.org/npm-conf/-/npm-conf-1.1.3.tgz",
      "integrity": "sha512-Yic4bZHJOt9RCFbRP3GgpqhScOY4HH3V2P8yBj6CeYq118Qr+BLXqT2JvpJ00mryLESpgOxf5XlFv4ZjXxLScw==",
      "requires": {
        "config-chain": "1.1.11",
        "pify": "3.0.0"
      }
    },
    "once": {
      "version": "1.4.0",
      "resolved": "https://registry.npmjs.org/once/-/once-1.4.0.tgz",
      "integrity": "sha1-WDsap3WWHUsROsF9nFC6753Xa9E=",
      "requires": {
        "wrappy": "1.0.2"
      }
    },
    "path-is-absolute": {
      "version": "1.0.1",
      "resolved": "https://registry.npmjs.org/path-is-absolute/-/path-is-absolute-1.0.1.tgz",
      "integrity": "sha1-F0uSaHNVNP+8es5r9TpanhtcX18="
    },
    "pify": {
      "version": "3.0.0",
      "resolved": "https://registry.npmjs.org/pify/-/pify-3.0.0.tgz",
      "integrity": "sha1-5aSs0sEB/fPZpNB/DbxNtJ3SgXY="
    },
    "prepend-http": {
      "version": "1.0.4",
      "resolved": "https://registry.npmjs.org/prepend-http/-/prepend-http-1.0.4.tgz",
      "integrity": "sha1-1PRWKwzjaW5BrFLQ4ALlemNdxtw="
    },
    "proto-list": {
      "version": "1.2.4",
      "resolved": "https://registry.npmjs.org/proto-list/-/proto-list-1.2.4.tgz",
      "integrity": "sha1-IS1b/hMYMGpCD2QCuOJv85ZHqEk="
    },
    "punycode": {
      "version": "1.3.2",
      "resolved": "https://registry.npmjs.org/punycode/-/punycode-1.3.2.tgz",
      "integrity": "sha1-llOgNvt8HuQjQvIyXM7v6jkmxI0=",
      "dev": true
    },
    "querystring": {
      "version": "0.2.0",
      "resolved": "https://registry.npmjs.org/querystring/-/querystring-0.2.0.tgz",
      "integrity": "sha1-sgmEkgO7Jd+CDadW50cAWHhSFiA=",
      "dev": true
    },
    "rimraf": {
      "version": "2.6.2",
      "resolved": "https://registry.npmjs.org/rimraf/-/rimraf-2.6.2.tgz",
      "integrity": "sha512-lreewLK/BlghmxtfH36YYVg1i8IAce4TI7oao75I1g245+6BctqTVQiBP3YUJ9C6DQOXJmkYR9X9fCLtCOJc5w==",
      "requires": {
        "glob": "7.1.2"
      }
    },
    "safe-buffer": {
      "version": "5.1.2",
      "resolved": "https://registry.npmjs.org/safe-buffer/-/safe-buffer-5.1.2.tgz",
      "integrity": "sha512-Gd2UZBJDkXlY7GbJxfsE8/nvKkUEU1G38c1siN6QP6a9PT9MmHB8GnpscSmMJSoF8LOIrt8ud/wPtojys4G6+g=="
    },
    "sax": {
      "version": "1.2.1",
      "resolved": "https://registry.npmjs.org/sax/-/sax-1.2.1.tgz",
      "integrity": "sha1-e45lYZCyKOgaZq6nSEgNgozS03o=",
      "dev": true
    },
    "semver": {
      "version": "5.5.0",
      "resolved": "https://registry.npmjs.org/semver/-/semver-5.5.0.tgz",
      "integrity": "sha512-4SJ3dm0WAwWy/NVeioZh5AntkdJoWKxHxcmyP622fOkgHa4z3R0TdBJICINyaSDE6uNwVc8gZr+ZinwZAH4xIA=="
    },
    "sharp": {
      "version": "0.17.3",
      "resolved": "https://registry.npmjs.org/sharp/-/sharp-0.17.3.tgz",
      "integrity": "sha1-SEzSpwyQA3CUjcxD4WX3gwa/9Io=",
      "requires": {
        "caw": "2.0.1",
        "color": "1.0.3",
        "got": "6.7.1",
        "nan": "2.10.0",
        "semver": "5.5.0",
        "tar": "2.2.1"
      }
    },
    "simple-swizzle": {
      "version": "0.2.2",
      "resolved": "https://registry.npmjs.org/simple-swizzle/-/simple-swizzle-0.2.2.tgz",
      "integrity": "sha1-pNprY1/8zMoz9w0Xy5JZLeleVXo=",
      "requires": {
        "is-arrayish": "0.3.2"
      }
    },
    "tar": {
      "version": "2.2.1",
      "resolved": "https://registry.npmjs.org/tar/-/tar-2.2.1.tgz",
      "integrity": "sha1-jk0qJWwOIYXGsYrWlK7JaLg8sdE=",
      "requires": {
        "block-stream": "0.0.9",
        "fstream": "1.0.11",
        "inherits": "2.0.3"
      }
    },
    "timed-out": {
      "version": "4.0.1",
      "resolved": "https://registry.npmjs.org/timed-out/-/timed-out-4.0.1.tgz",
      "integrity": "sha1-8y6srFoXW+ol1/q1Zas+2HQe9W8="
    },
    "tunnel-agent": {
      "version": "0.6.0",
      "resolved": "https://registry.npmjs.org/tunnel-agent/-/tunnel-agent-0.6.0.tgz",
      "integrity": "sha1-J6XeoGs2sEoKmWZ3SykIaPD8QP0=",
      "requires": {
        "safe-buffer": "5.1.2"
      }
    },
    "unzip-response": {
      "version": "2.0.1",
      "resolved": "https://registry.npmjs.org/unzip-response/-/unzip-response-2.0.1.tgz",
      "integrity": "sha1-0vD3N9FrBhXnKmk17QQhRXLVb5c="
    },
    "url": {
      "version": "0.10.3",
      "resolved": "https://registry.npmjs.org/url/-/url-0.10.3.tgz",
      "integrity": "sha1-Ah5NnHcF8hu/N9A861h2dAJ3TGQ=",
      "dev": true,
      "requires": {
        "punycode": "1.3.2",
        "querystring": "0.2.0"
      }
    },
    "url-parse-lax": {
      "version": "1.0.0",
      "resolved": "https://registry.npmjs.org/url-parse-lax/-/url-parse-lax-1.0.0.tgz",
      "integrity": "sha1-evjzA2Rem9eaJy56FKxovAYJ2nM=",
      "requires": {
        "prepend-http": "1.0.4"
      }
    },
    "url-to-options": {
      "version": "1.0.1",
      "resolved": "https://registry.npmjs.org/url-to-options/-/url-to-options-1.0.1.tgz",
      "integrity": "sha1-FQWgOiiaSMvXpDTvuu7FBV9WM6k="
    },
    "uuid": {
      "version": "3.1.0",
      "resolved": "https://registry.npmjs.org/uuid/-/uuid-3.1.0.tgz",
      "integrity": "sha512-DIWtzUkw04M4k3bf1IcpS2tngXEL26YUD2M0tMDUpnUrz2hgzUBlD55a4FjdLGPvfHxS6uluGWvaVEqgBcVa+g==",
      "dev": true
    },
    "wrappy": {
      "version": "1.0.2",
      "resolved": "https://registry.npmjs.org/wrappy/-/wrappy-1.0.2.tgz",
      "integrity": "sha1-tSQ9jz7BqjXxNkYFvA0QNuMKtp8="
    },
    "xml2js": {
      "version": "0.4.17",
      "resolved": "https://registry.npmjs.org/xml2js/-/xml2js-0.4.17.tgz",
      "integrity": "sha1-F76T6q4/O3eTWceVtBlwWogX6Gg=",
      "dev": true,
      "requires": {
        "sax": "1.2.1",
        "xmlbuilder": "4.2.1"
      }
    },
    "xmlbuilder": {
      "version": "4.2.1",
      "resolved": "https://registry.npmjs.org/xmlbuilder/-/xmlbuilder-4.2.1.tgz",
      "integrity": "sha1-qlijBBoGb5DqoWwvU4n/GfP0YaU=",
      "dev": true,
      "requires": {
        "lodash": "4.17.10"
      }
    }
  }
}
